module adder(intput a,
    input b,
    output sum);
endmodule